** PMOS transfer characteristics
Vg 1 0 dc -2v
Vd 3 0 dc -2.5v
V1 3 2 dc 0v
.model pmod pmos level = 54 version = 4.7
M1 0 1 2 2 pmod w = 100u l = 10u
.dc Vd 0 -2.5 -0.1 Vg 0 -2.0 -0.1
.control
run
plot i(V1)
.endc
.end 