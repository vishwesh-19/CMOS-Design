** 3 Input NOR Gate
Vd 5 0 dc 5V
V1 1 0 pulse(0 5 0 0 0 10m 20m)
V2 2 0 pulse(0 5 0 0 0 5m 20m)
V3 3 0 pulse(0 5 0 0 0 15m 20m)
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
m1a 4 1 0 0 nmod w=100u l=10u
m2b 4 2 0 0 nmod w=100u l=10u
m2c 4 3 0 0 nmod w=100u l=10u
m2a 6 1 5 5 pmod w=100u l=10u
m2b 7 2 6 5 pmod w=100u l=10u
m2c 4 3 7 5 pmod w=100u l=10u
.tran 0.1m 100m
.control
run
plot V(1) V(2) V(3) 
plot V(4)
.endc
.end