** CMOS Inverter Characteristics
Vg 1 0 5.0
Vd 3 0 dc 5v
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
m1 2 1 0 0 nmod w=100u l=10u
m2 2 1 3 3 pmod w=100u l=10u
.dc Vg 0.0 5.0 0.1 
.control
run
plot V(1) V(2)
.endc
.end